package instr_agent_pkg;
`include "uvm_macros.svh"
import uvm_pkg::*;
import tb_top_pkg::*;

`include "instr_packet.sv"
`include "instr_driver.sv"
`include "instr_monitor.sv"
`include "instr_seqr.sv"
`include "instr_agent_cfg.sv" 
`include "instr_agent.sv" 

endpackage
