// ***************************************************
//    TB_TOP package
// ***************************************************


package tb_top_pkg;
`include "uvm_macros.svh"
import uvm_pkg::*;

endpackage
