package tb_scoreboard_pkg;

`include "uvm_macros.svh"
import uvm_pkg::*;
import instr_agent_pkg::*;
import load_agent_pkg::*;

`include "tb_scoreboard.sv"

endpackage
