package load_req_resp_agent_pkg;

`include "uvm_macros.svh"
import uvm_pkg::*;
import tb_top_pkg::*;

`include "load_req_resp_packet.sv"
`include "load_req_resp_monitor.sv"
`include "load_req_resp_driver.sv"
`include "load_req_resp_sequencer.sv"
`include "load_req_resp_agent_config.sv"
`include "load_req_resp_agent.sv"
`include "load_req_resp_sequence.sv"
endpackage
