package tb_test_pkg;

`include "uvm_macros.svh"
import uvm_pkg::*;
import tb_top_pkg::*;
import tb_env_pkg::*;

`include "test_base.sv"

endpackage
