`ifndef DEFINES_SVH
`define DEFINES_SVH

`define FIFO_DEPTH 4
`define REG_WIDTH  5
`define OP_WIDTH   5

typedef enum bit { 
   UVM_PASSIVE=0, 
   UVM_ACTIVE=1
} uvm_active_passive_enum;

`endif
