package load_agent_pkg;

`include "uvm_macros.svh"
import uvm_pkg::*;
import tb_top_pkg::*;

`include "load_packet.sv"
`include "load_monitor.sv"
`include "load_slave_driver.sv"
`include "load_sequencer.sv"
`include "load_sequence.sv"
`include "load_agent_cfg.sv"
`include "load_agent.sv"


endpackage