// ENV package.. 
//
package tb_env_pkg; 
`include "uvm_macros.svh"
import uvm_pkg::*;
import instr_agent_pkg::*;
import load_agent_pkg::*;
import tb_sequences_pkg::*;
import tb_scoreboard_pkg::*;

`include "tb_env.sv"

endpackage
